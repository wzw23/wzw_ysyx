	// verilator_coverage annotation
%000067	module Alu(input [63:0]a, input [63:0]b,output [63:0]out);
%000041	verilator_coverage: (next point on previous line)

%000068	verilator_coverage: (next point on previous line)

	    assign out=a+b;
	endmodule
	
