	// verilator_coverage annotation
	// 带默认值的选择器模板
	module MuxKeyWithDefault #(NR_KEY = 2, KEY_LEN = 1, DATA_LEN = 1) (
%000041	  output [DATA_LEN-1:0] out,
%000004	  input [KEY_LEN-1:0] key,
%000000	  input [DATA_LEN-1:0] default_out,
	  input [NR_KEY*(KEY_LEN + DATA_LEN)-1:0] lut
	);
	  MuxKeyInternal #(NR_KEY, KEY_LEN, DATA_LEN, 1) i0 (out, key, default_out, lut);
	endmodule
	
